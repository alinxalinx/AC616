//===========================================================================
// Module name: io_test.v
// ����: 0.5������IO��ƽ��0.5������IO��ƽ
//===========================================================================
`timescale 1ns / 1ps

module io_test (
                  clk,           // ������������ʱ��: 50Mhz
                  rst_n,         // �����������븴λ����
                  j3_io,         // ���ڿ��ƿ�������J3�������ϵ�IO
                  j4_io,         // ���ڿ��ƿ�������J4�������ϵ�IO
                  j6_io,         // ���ڿ��ƿ�������J6�������ϵ�IO
                  j7_io         // ���ڿ��ƿ�������J7�������ϵ�IO						
             );
             
//===========================================================================
// PORT declarations
//===========================================================================
input clk;
input rst_n;
output [33:0] j3_io;
output [33:0] j4_io;
output [33:0] j6_io;
output [33:0] j7_io;

//�Ĵ�������
reg [31:0] timer;    
              
reg [33:0] j3_io_reg;
reg [33:0] j4_io_reg;
reg [33:0] j6_io_reg;
reg [33:0] j7_io_reg;

assign j3_io=j3_io_reg;
assign j4_io=j4_io_reg;
assign j6_io=j6_io_reg;
assign j7_io=j7_io_reg;
//===========================================================================
// ����������:ѭ������0~4��
//===========================================================================
  always @(posedge clk or negedge rst_n)    //���ʱ�ӵ������غ͸�λ���½���
    begin
      if (~rst_n)                           //��λ�źŵ���Ч
          timer <= 0;                       //����������
      else if (timer == 32'd24_999_999)    //������ʹ�õľ���Ϊ50MHz��0.5�����(50M*0.5-1=24_999_999)
          timer <= 0;                       //�������Ƶ�4�룬����������
      else
		    timer <= timer + 1'b1;            //��������1
    end

//===========================================================================
// LED�ƿ���
//===========================================================================
  always @(posedge clk or negedge rst_n)   //���ʱ�ӵ������غ͸�λ���½���
    begin
      if (~rst_n) begin                    //��λ�źŵ���Ч
		   j3_io_reg<=0;                     //IOȫΪ�͵�ƽ
		   j4_io_reg<=0;                     //IOȫΪ�͵�ƽ
		   j6_io_reg<=0;                     //IOȫΪ�͵�ƽ  
		   j7_io_reg<=0;                     //IOȫΪ�͵�ƽ 
      end			
      else if (timer == 32'd24_999_999) begin    //�������Ƶ�1�룬
		   j3_io_reg<=~j3_io_reg;                  //IO��ƽ��ת
		   j4_io_reg<=~j4_io_reg;                  //IO��ƽ��ת
		   j6_io_reg<=~j6_io_reg;                  //IO��ƽ��ת 
		   j7_io_reg<=~j7_io_reg;                  //IO��ƽ��ת 
		end   
    end
    
endmodule

