//===========================================================================
// Module name: led_test.v
// ����: ÿ��1�����ε����������ϵ�LED0~LED4
//===========================================================================
`timescale 1ns / 1ps

module led_test (
                  clk,           // ������������ʱ��: 50Mhz
                  rst_n,         // �����������븴λ����
                  led            // ���LED��,���ڿ��ƿ��������ĸ�LED(LED1~LED4)
             );
             
//===========================================================================
// PORT declarations
//===========================================================================
input clk;
input rst_n;
output [3:0] led;

//�Ĵ�������
reg [31:0] timer;                  
reg [3:0] led;


//===========================================================================
// ����������:ѭ������0~4��
//===========================================================================
  always @(posedge clk or negedge rst_n)    //���ʱ�ӵ������غ͸�λ���½���
    begin
      if (~rst_n)                           //��λ�źŵ���Ч
          timer <= 0;                       //����������
      else if (timer == 32'd199_999_999)    //������ʹ�õľ���Ϊ50MHz��4�����(50M*4-1=199_999_999)
          timer <= 0;                       //�������Ƶ�4�룬����������
      else
		    timer <= timer + 1'b1;            //��������1
    end

//===========================================================================
// LED�ƿ���
//===========================================================================
  always @(posedge clk or negedge rst_n)   //���ʱ�ӵ������غ͸�λ���½���
    begin
      if (~rst_n)                          //��λ�źŵ���Ч
          led <= 4'b1111;                  //LED�����ȫΪ�ߣ��ĸ�LED����           
      else if (timer == 32'd49_999_999)    //�������Ƶ�1�룬
          led <= 4'b1110;                  //LED1����
      else if (timer == 32'd99_999_999)    //�������Ƶ�2�룬
          led <= 4'b1101;                  //LED2����
      else if (timer == 32'd149_999_999)   //�������Ƶ�3�룬
          led <= 4'b1011;                  //LED3����                           
      else if (timer == 32'd199_999_999)   //�������Ƶ�4�룬
          led <= 4'b0111;                  //LED4����        
    end
    
endmodule

